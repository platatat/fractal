module DE1_SoC_Computer (
	////////////////////////////////////
	// FPGA Pins
	////////////////////////////////////

	// Clock pins
	CLOCK_50,
	CLOCK2_50,
	CLOCK3_50,
	CLOCK4_50,

	// ADC
	ADC_CS_N,
	ADC_DIN,
	ADC_DOUT,
	ADC_SCLK,

	// Audio
	AUD_ADCDAT,
	AUD_ADCLRCK,
	AUD_BCLK,
	AUD_DACDAT,
	AUD_DACLRCK,
	AUD_XCK,

	// SDRAM
	DRAM_ADDR,
	DRAM_BA,
	DRAM_CAS_N,
	DRAM_CKE,
	DRAM_CLK,
	DRAM_CS_N,
	DRAM_DQ,
	DRAM_LDQM,
	DRAM_RAS_N,
	DRAM_UDQM,
	DRAM_WE_N,

	// I2C Bus for Configuration of the Audio and Video-In Chips
	FPGA_I2C_SCLK,
	FPGA_I2C_SDAT,

	// 40-Pin Headers
	GPIO_0,
	GPIO_1,
	
	// Seven Segment Displays
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,

	// IR
	IRDA_RXD,
	IRDA_TXD,

	// Pushbuttons
	KEY,

	// LEDs
	LEDR,

	// PS2 Ports
	PS2_CLK,
	PS2_DAT,
	
	PS2_CLK2,
	PS2_DAT2,

	// Slider Switches
	SW,

	// Video-In
	TD_CLK27,
	TD_DATA,
	TD_HS,
	TD_RESET_N,
	TD_VS,

	// VGA
	VGA_B,
	VGA_BLANK_N,
	VGA_CLK,
	VGA_G,
	VGA_HS,
	VGA_R,
	VGA_SYNC_N,
	VGA_VS,

	////////////////////////////////////
	// HPS Pins
	////////////////////////////////////
	
	// DDR3 SDRAM
	HPS_DDR3_ADDR,
	HPS_DDR3_BA,
	HPS_DDR3_CAS_N,
	HPS_DDR3_CKE,
	HPS_DDR3_CK_N,
	HPS_DDR3_CK_P,
	HPS_DDR3_CS_N,
	HPS_DDR3_DM,
	HPS_DDR3_DQ,
	HPS_DDR3_DQS_N,
	HPS_DDR3_DQS_P,
	HPS_DDR3_ODT,
	HPS_DDR3_RAS_N,
	HPS_DDR3_RESET_N,
	HPS_DDR3_RZQ,
	HPS_DDR3_WE_N,

	// Ethernet
	HPS_ENET_GTX_CLK,
	HPS_ENET_INT_N,
	HPS_ENET_MDC,
	HPS_ENET_MDIO,
	HPS_ENET_RX_CLK,
	HPS_ENET_RX_DATA,
	HPS_ENET_RX_DV,
	HPS_ENET_TX_DATA,
	HPS_ENET_TX_EN,

	// Flash
	HPS_FLASH_DATA,
	HPS_FLASH_DCLK,
	HPS_FLASH_NCSO,

	// Accelerometer
	HPS_GSENSOR_INT,
		
	// General Purpose I/O
	HPS_GPIO,
		
	// I2C
	HPS_I2C_CONTROL,
	HPS_I2C1_SCLK,
	HPS_I2C1_SDAT,
	HPS_I2C2_SCLK,
	HPS_I2C2_SDAT,

	// Pushbutton
	HPS_KEY,

	// LED
	HPS_LED,
		
	// SD Card
	HPS_SD_CLK,
	HPS_SD_CMD,
	HPS_SD_DATA,

	// SPI
	HPS_SPIM_CLK,
	HPS_SPIM_MISO,
	HPS_SPIM_MOSI,
	HPS_SPIM_SS,

	// UART
	HPS_UART_RX,
	HPS_UART_TX,

	// USB
	HPS_CONV_USB_N,
	HPS_USB_CLKOUT,
	HPS_USB_DATA,
	HPS_USB_DIR,
	HPS_USB_NXT,
	HPS_USB_STP
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

////////////////////////////////////
// FPGA Pins
////////////////////////////////////

// Clock pins
input						CLOCK_50;
input						CLOCK2_50;
input						CLOCK3_50;
input						CLOCK4_50;

// ADC
inout						ADC_CS_N;
output					ADC_DIN;
input						ADC_DOUT;
output					ADC_SCLK;

// Audio
input						AUD_ADCDAT;
inout						AUD_ADCLRCK;
inout						AUD_BCLK;
output					AUD_DACDAT;
inout						AUD_DACLRCK;
output					AUD_XCK;

// SDRAM
output 		[12: 0]	DRAM_ADDR;
output		[ 1: 0]	DRAM_BA;
output					DRAM_CAS_N;
output					DRAM_CKE;
output					DRAM_CLK;
output					DRAM_CS_N;
inout			[15: 0]	DRAM_DQ;
output					DRAM_LDQM;
output					DRAM_RAS_N;
output					DRAM_UDQM;
output					DRAM_WE_N;

// I2C Bus for Configuration of the Audio and Video-In Chips
output					FPGA_I2C_SCLK;
inout						FPGA_I2C_SDAT;

// 40-pin headers
inout			[35: 0]	GPIO_0;
inout			[35: 0]	GPIO_1;

// Seven Segment Displays
output		[ 6: 0]	HEX0;
output		[ 6: 0]	HEX1;
output		[ 6: 0]	HEX2;
output		[ 6: 0]	HEX3;
output		[ 6: 0]	HEX4;
output		[ 6: 0]	HEX5;

// IR
input						IRDA_RXD;
output					IRDA_TXD;

// Pushbuttons
input			[ 3: 0]	KEY;

// LEDs
output		[ 9: 0]	LEDR;

// PS2 Ports
inout						PS2_CLK;
inout						PS2_DAT;

inout						PS2_CLK2;
inout						PS2_DAT2;

// Slider Switches
input			[ 9: 0]	SW;

// Video-In
input						TD_CLK27;
input			[ 7: 0]	TD_DATA;
input						TD_HS;
output					TD_RESET_N;
input						TD_VS;

// VGA
output		[ 7: 0]	VGA_B;
output					VGA_BLANK_N;
output					VGA_CLK;
output		[ 7: 0]	VGA_G;
output					VGA_HS;
output		[ 7: 0]	VGA_R;
output					VGA_SYNC_N;
output					VGA_VS;



////////////////////////////////////
// HPS Pins
////////////////////////////////////
	
// DDR3 SDRAM
output		[14: 0]	HPS_DDR3_ADDR;
output		[ 2: 0]  HPS_DDR3_BA;
output					HPS_DDR3_CAS_N;
output					HPS_DDR3_CKE;
output					HPS_DDR3_CK_N;
output					HPS_DDR3_CK_P;
output					HPS_DDR3_CS_N;
output		[ 3: 0]	HPS_DDR3_DM;
inout			[31: 0]	HPS_DDR3_DQ;
inout			[ 3: 0]	HPS_DDR3_DQS_N;
inout			[ 3: 0]	HPS_DDR3_DQS_P;
output					HPS_DDR3_ODT;
output					HPS_DDR3_RAS_N;
output					HPS_DDR3_RESET_N;
input						HPS_DDR3_RZQ;
output					HPS_DDR3_WE_N;

// Ethernet
output					HPS_ENET_GTX_CLK;
inout						HPS_ENET_INT_N;
output					HPS_ENET_MDC;
inout						HPS_ENET_MDIO;
input						HPS_ENET_RX_CLK;
input			[ 3: 0]	HPS_ENET_RX_DATA;
input						HPS_ENET_RX_DV;
output		[ 3: 0]	HPS_ENET_TX_DATA;
output					HPS_ENET_TX_EN;

// Flash
inout			[ 3: 0]	HPS_FLASH_DATA;
output					HPS_FLASH_DCLK;
output					HPS_FLASH_NCSO;

// Accelerometer
inout						HPS_GSENSOR_INT;

// General Purpose I/O
inout			[ 1: 0]	HPS_GPIO;

// I2C
inout						HPS_I2C_CONTROL;
inout						HPS_I2C1_SCLK;
inout						HPS_I2C1_SDAT;
inout						HPS_I2C2_SCLK;
inout						HPS_I2C2_SDAT;

// Pushbutton
inout						HPS_KEY;

// LED
inout						HPS_LED;

// SD Card
output					HPS_SD_CLK;
inout						HPS_SD_CMD;
inout			[ 3: 0]	HPS_SD_DATA;

// SPI
output					HPS_SPIM_CLK;
input						HPS_SPIM_MISO;
output					HPS_SPIM_MOSI;
inout						HPS_SPIM_SS;

// UART
input						HPS_UART_RX;
output					HPS_UART_TX;

// USB
inout						HPS_CONV_USB_N;
input						HPS_USB_CLKOUT;
inout			[ 7: 0]	HPS_USB_DATA;
input						HPS_USB_DIR;
input						HPS_USB_NXT;
output					HPS_USB_STP;

//=======================================================
//  REG/WIRE declarations
//=======================================================

wire			[23: 0]	hex5_hex0;
//wire			[15: 0]	hex5_hex4;

//assign HEX0 = ~hex3_hex0[ 6: 0]; // hex3_hex0[ 6: 0]; 
//assign HEX1 = ~hex3_hex0[14: 8];
//assign HEX2 = ~hex3_hex0[22:16];
//assign HEX3 = ~hex3_hex0[30:24];
//assign HEX4 = 7'b1111111;
//assign HEX5 = 7'b1111111;

HexDigit Digit0(HEX0, hex5_hex0[3:0]);
HexDigit Digit1(HEX1, hex5_hex0[7:4]);
HexDigit Digit2(HEX2, hex5_hex0[11:8]);
HexDigit Digit3(HEX3, hex5_hex0[15:12]);
HexDigit Digit4(HEX4, hex5_hex0[19:16]);
HexDigit Digit5(HEX5, hex5_hex0[23:20]);

//=======================================================
// OLD Solvers and VGA logic
//=======================================================
wire reset_key;
assign reset_key = ~KEY[0];

// wire stream_ready;
// wire stream_start;
// wire stream_end;
// wire stream_valid;

// wire [15:0] stream_data;

// wire [5:0] solver_id;
// wire [18:0] solver_addr;

// localparam NUM_SOLVERS = 29;

// pixel_iterator #(NUM_SOLVERS, 640, 480) pixel_it (
//     .clock(CLOCK_50),
//     .reset(reset_key),
//     .en(stream_ready),

//     .solver_id(solver_id),
//     .solver_addr(solver_addr),

//     .start_stream(stream_start),
//     .end_stream(stream_end),
//     .valid_stream(stream_valid)
// );

reg stream_start_delay [2:1];
reg stream_end_delay [2:1];
reg stream_valid_delay [2:1];

// always @(posedge CLOCK_50) begin
//     stream_start_delay[1] <= stream_start;
//     stream_end_delay[1] <= stream_end;
//     stream_valid_delay[1] <= stream_valid;

//     stream_start_delay[2] <= stream_start_delay[1];
//     stream_end_delay[2] <= stream_end_delay[1];
//     stream_valid_delay[2] <= stream_valid_delay[1];
// end

// wire [31:0] solve_time;
// reg signed [3:0] solver_data_out;

// wire signed [26:0] x_min, y_min;
// wire signed [26:0] dx, dy;

// wire [9:0] solver_iterations;
// wire solver_hps_reset;
// wire solver_done;
// wire solver_clock;

// multi_solver #(NUM_SOLVERS) solver (
//     .clock(solver_clock),
//     .reset(reset_key | solver_hps_reset),

//     .min_x(x_min),
//     .min_y(y_min),
//     .dx(dx),
//     .dy(dy),
//     .iterations(solver_iterations),

//     .rd_clock(CLOCK_50),
//     .rd_solver_id(solver_id),
//     .rd_addr(solver_addr),
//     .rd_data_out(solver_data_out),

//     .solve_time(solve_time),
//     .done(solver_done)
// );

// assign stream_data = {5'b0, solver_data_out, 7'b0};

// assign stream_data = 
// 		solver_data_out == 4'b0000 ? 16'b00000_000000_00000 :
// 		solver_data_out == 4'b0001 ? 16'b00000_001000_00000 :
// 		solver_data_out == 4'b0010 ? 16'b00000_010000_00000 :
// 		solver_data_out == 4'b0011 ? 16'b00000_011000_00000 :
// 		solver_data_out == 4'b0100 ? 16'b00000_100000_00000 :
// 		solver_data_out == 4'b0101 ? 16'b00000_101000_00000 :
// 		solver_data_out == 4'b0110 ? 16'b00000_110000_00000 :
// 		solver_data_out == 4'b0111 ? 16'b00000_111000_01000 :
// 		solver_data_out == 4'b1000 ? 16'b00000_111000_10000 :
// 		solver_data_out == 4'b1001 ? 16'b00000_110000_11000 :
// 		solver_data_out == 4'b1010 ? 16'b00000_101000_11000 :
// 		solver_data_out == 4'b1011 ? 16'b00000_100000_11000 :
// 		solver_data_out == 4'b1100 ? 16'b00000_011000_11000 :
// 		solver_data_out == 4'b1101 ? 16'b00000_010000_11000 :
// 		solver_data_out == 4'b1110 ? 16'b00000_001000_11000 :
// 		solver_data_out == 4'b1111 ? 16'b00000_000000_11000 :
// 									 16'b11111_000000_00000;

// assign hex5_hex0 = solve_time[23:0];
// assign LEDR[7:0] = solve_time[31:24];

//=======================================================
// NEW Solvers and VGA logic
//=======================================================

localparam NUM_SOLVERS 			= 2;
localparam TILE_WIDTH_BITS      = 6;
localparam LIMB_INDEX_BITS 		= 6;
localparam LIMB_SIZE_BITS 		= 27;
localparam DIVERGENCE_RADIUS 	= 4;

wire [31:0] fifo_raw_data;
wire        fifo_valid;
wire        fifo_ready;
wire        fifo_startofpacket;
wire        fifo_endofpacket;

/*
wire [2:0] 	fifo_data_type;
wire [31:0] fifo_decoded_data;

hps_fifo_decoder hps_fifo_decoder (
	.raw_data 		(fifo_raw_data),
	.data_type 		(fifo_data_type),
	.decoded_data 	(fifo_decoded_data)
);

solver_manager #(
	NUM_SOLVERS,
	LIMB_INDEX_BITS,
	LIMB_SIZE_BITS,
	DIVERGENCE_RADIUS
) solver_manager (
	.clock 			(CLOCK_50),
	.reset 			(~KEY[0]),
	.fifo_valid 	(fifo_valid),
	.fifo_data_type (fifo_data_type),
	.fifo_data 		(fifo_decoded_data),
	.fifo_ready     (fifo_ready)
);
*/

/*
wire [15:0] write_out_data;
wire [31:0] write_out_addr;
wire write_out_ready;
wire write_out_valid;

tile_solver_legit #(
    TILE_WIDTH_BITS,
	LIMB_INDEX_BITS,
	LIMB_SIZE_BITS,
	DIVERGENCE_RADIUS
) tile_solver(
    .clock(CLOCK_50),
    .reset(reset_key),

    .in_data(fifo_raw_data),
    .in_valid(fifo_valid),
    .in_ready(fifo_ready),
    .in_end_of_stream(fifo_endofpacket),

    .out_addr(write_out_addr),
    .out_data(write_out_data),
    .out_valid(write_out_valid),
    .out_ready(write_out_ready)
);

reg [1:0] state;
reg [31:0] write_addr;
reg [15:0] write_data;
wire write_en;
wire ack;

always @(posedge CLOCK_50) begin
    if (reset_key) begin
        state <= 0;
        write_addr <= 0;
        write_data <= 0;
    end else if (state == 0) begin
        // Wait for data
        if (write_out_valid) begin
            state <= 1;
            write_data <= write_out_data;
            write_addr <= write_out_addr;
        end else begin
            state <= 0;
        end
    end else if (state == 1) begin
        // Wait for ack
        if (ack) begin
            state <= 0;
        end else begin
            state <= 1;
        end
    end
end

assign write_en = (state == 1);
assign write_out_ready = (state == 0);
*/

wire [31:0] in_data;
wire        in_valid;
wire        in_end_of_stream;
wire        in_ready;

wire [15:0] out_data;
wire [31:0] out_addr;
wire        out_write_en;
wire        out_ack;

multi_tile_solver #(
    NUM_SOLVERS,
    TILE_WIDTH_BITS,
    LIMB_INDEX_BITS,
    LIMB_SIZE_BITS,
    DIVERGENCE_RADIUS
) (
    .clock(CLOCK_50),
    .reset(reset_key),

    .in_data(in_data),
    .in_valid(in_valid),
    .in_end_of_stream(in_end_of_stream),
    .in_ready(in_ready),

    .out_data(out_data),
    .out_addr(out_addr),
    .out_write_en(out_write_en),
    .out_ack(out_ack)
);

//=======================================================
//  Structural coding
//=======================================================
// From Qsys

Computer_System The_System (
	////////////////////////////////////
	// FPGA Side
	////////////////////////////////////

	// Global signals
	.system_pll_ref_clk_clk					(CLOCK_50),
	.system_pll_ref_reset_reset			(1'b0),
	
	// SDRAM
	.sdram_clk_clk								(DRAM_CLK),
	.sdram_addr									(DRAM_ADDR),
	.sdram_ba									(DRAM_BA),
	.sdram_cas_n								(DRAM_CAS_N),
	.sdram_cke									(DRAM_CKE),
	.sdram_cs_n									(DRAM_CS_N),
	.sdram_dq									(DRAM_DQ),
	.sdram_dqm									({DRAM_UDQM,DRAM_LDQM}),
	.sdram_ras_n								(DRAM_RAS_N),
	.sdram_we_n									(DRAM_WE_N),

	////////////////////////////////////
	// HPS Side
	////////////////////////////////////
	// DDR3 SDRAM
	.memory_mem_a			(HPS_DDR3_ADDR),
	.memory_mem_ba			(HPS_DDR3_BA),
	.memory_mem_ck			(HPS_DDR3_CK_P),
	.memory_mem_ck_n		(HPS_DDR3_CK_N),
	.memory_mem_cke		(HPS_DDR3_CKE),
	.memory_mem_cs_n		(HPS_DDR3_CS_N),
	.memory_mem_ras_n		(HPS_DDR3_RAS_N),
	.memory_mem_cas_n		(HPS_DDR3_CAS_N),
	.memory_mem_we_n		(HPS_DDR3_WE_N),
	.memory_mem_reset_n	(HPS_DDR3_RESET_N),
	.memory_mem_dq			(HPS_DDR3_DQ),
	.memory_mem_dqs		(HPS_DDR3_DQS_P),
	.memory_mem_dqs_n		(HPS_DDR3_DQS_N),
	.memory_mem_odt		(HPS_DDR3_ODT),
	.memory_mem_dm			(HPS_DDR3_DM),
	.memory_oct_rzqin		(HPS_DDR3_RZQ),
		  
	// Ethernet
	.hps_io_hps_io_gpio_inst_GPIO35	(HPS_ENET_INT_N),
	.hps_io_hps_io_emac1_inst_TX_CLK	(HPS_ENET_GTX_CLK),
	.hps_io_hps_io_emac1_inst_TXD0	(HPS_ENET_TX_DATA[0]),
	.hps_io_hps_io_emac1_inst_TXD1	(HPS_ENET_TX_DATA[1]),
	.hps_io_hps_io_emac1_inst_TXD2	(HPS_ENET_TX_DATA[2]),
	.hps_io_hps_io_emac1_inst_TXD3	(HPS_ENET_TX_DATA[3]),
	.hps_io_hps_io_emac1_inst_RXD0	(HPS_ENET_RX_DATA[0]),
	.hps_io_hps_io_emac1_inst_MDIO	(HPS_ENET_MDIO),
	.hps_io_hps_io_emac1_inst_MDC		(HPS_ENET_MDC),
	.hps_io_hps_io_emac1_inst_RX_CTL	(HPS_ENET_RX_DV),
	.hps_io_hps_io_emac1_inst_TX_CTL	(HPS_ENET_TX_EN),
	.hps_io_hps_io_emac1_inst_RX_CLK	(HPS_ENET_RX_CLK),
	.hps_io_hps_io_emac1_inst_RXD1	(HPS_ENET_RX_DATA[1]),
	.hps_io_hps_io_emac1_inst_RXD2	(HPS_ENET_RX_DATA[2]),
	.hps_io_hps_io_emac1_inst_RXD3	(HPS_ENET_RX_DATA[3]),

	// Flash
	.hps_io_hps_io_qspi_inst_IO0	(HPS_FLASH_DATA[0]),
	.hps_io_hps_io_qspi_inst_IO1	(HPS_FLASH_DATA[1]),
	.hps_io_hps_io_qspi_inst_IO2	(HPS_FLASH_DATA[2]),
	.hps_io_hps_io_qspi_inst_IO3	(HPS_FLASH_DATA[3]),
	.hps_io_hps_io_qspi_inst_SS0	(HPS_FLASH_NCSO),
	.hps_io_hps_io_qspi_inst_CLK	(HPS_FLASH_DCLK),

	// Accelerometer
	.hps_io_hps_io_gpio_inst_GPIO61	(HPS_GSENSOR_INT),

	//.adc_sclk                        (ADC_SCLK),
	//.adc_cs_n                        (ADC_CS_N),
	//.adc_dout                        (ADC_DOUT),
	//.adc_din                         (ADC_DIN),

	// General Purpose I/O
	.hps_io_hps_io_gpio_inst_GPIO40	(HPS_GPIO[0]),
	.hps_io_hps_io_gpio_inst_GPIO41	(HPS_GPIO[1]),

	// I2C
	.hps_io_hps_io_gpio_inst_GPIO48	(HPS_I2C_CONTROL),
	.hps_io_hps_io_i2c0_inst_SDA		(HPS_I2C1_SDAT),
	.hps_io_hps_io_i2c0_inst_SCL		(HPS_I2C1_SCLK),
	.hps_io_hps_io_i2c1_inst_SDA		(HPS_I2C2_SDAT),
	.hps_io_hps_io_i2c1_inst_SCL		(HPS_I2C2_SCLK),

	// Pushbutton
	.hps_io_hps_io_gpio_inst_GPIO54	(HPS_KEY),

	// LED
	.hps_io_hps_io_gpio_inst_GPIO53	(HPS_LED),

	// SD Card
	.hps_io_hps_io_sdio_inst_CMD	(HPS_SD_CMD),
	.hps_io_hps_io_sdio_inst_D0	(HPS_SD_DATA[0]),
	.hps_io_hps_io_sdio_inst_D1	(HPS_SD_DATA[1]),
	.hps_io_hps_io_sdio_inst_CLK	(HPS_SD_CLK),
	.hps_io_hps_io_sdio_inst_D2	(HPS_SD_DATA[2]),
	.hps_io_hps_io_sdio_inst_D3	(HPS_SD_DATA[3]),

	// SPI
	.hps_io_hps_io_spim1_inst_CLK		(HPS_SPIM_CLK),
	.hps_io_hps_io_spim1_inst_MOSI	(HPS_SPIM_MOSI),
	.hps_io_hps_io_spim1_inst_MISO	(HPS_SPIM_MISO),
	.hps_io_hps_io_spim1_inst_SS0		(HPS_SPIM_SS),

	// UART
	.hps_io_hps_io_uart0_inst_RX	(HPS_UART_RX),
	.hps_io_hps_io_uart0_inst_TX	(HPS_UART_TX),

	// USB
	.hps_io_hps_io_gpio_inst_GPIO09	(HPS_CONV_USB_N),
	.hps_io_hps_io_usb1_inst_D0		(HPS_USB_DATA[0]),
	.hps_io_hps_io_usb1_inst_D1		(HPS_USB_DATA[1]),
	.hps_io_hps_io_usb1_inst_D2		(HPS_USB_DATA[2]),
	.hps_io_hps_io_usb1_inst_D3		(HPS_USB_DATA[3]),
	.hps_io_hps_io_usb1_inst_D4		(HPS_USB_DATA[4]),
	.hps_io_hps_io_usb1_inst_D5		(HPS_USB_DATA[5]),
	.hps_io_hps_io_usb1_inst_D6		(HPS_USB_DATA[6]),
	.hps_io_hps_io_usb1_inst_D7		(HPS_USB_DATA[7]),
	.hps_io_hps_io_usb1_inst_CLK		(HPS_USB_CLKOUT),
	.hps_io_hps_io_usb1_inst_STP		(HPS_USB_STP),
	.hps_io_hps_io_usb1_inst_DIR		(HPS_USB_DIR),
	.hps_io_hps_io_usb1_inst_NXT		(HPS_USB_NXT),

    .sdram_writer_address     (out_addr),
    .sdram_writer_byte_enable (2'b11),
    .sdram_writer_write       (out_write_en),
    .sdram_writer_write_data  (out_data),
    .sdram_writer_acknowledge (out_ack),
    //.sdram_writer_read        (),
    //.sdram_writer_read_data   (),

    .in_fifo_data  (in_data),
    .in_fifo_valid (in_valid),
    .in_fifo_ready (in_ready),
    .in_fifo_startofpacket (),
    .in_fifo_endofpacket   (in_end_of_stream),
);
endmodule // end top level
